/*
* LineBuf.sv
* Author: Aero2021
* Version: 2.0: 固定bram的深度    
*/

`timescale 1ns / 1ps

module LineBuf #(
    parameter DATA_WIDTH = 8,
    parameter LATENCY = 0
) (
    input   clk,
    input   rst_n,
    input   in_valid,
    input  [DATA_WIDTH-1:0] data_in,
    output [DATA_WIDTH-1:0] data_out
);
    localparam ADDR_WIDTH = $clog2(LATENCY);
    localparam BRAM_DEPTH = 8192;

    initial begin
        if (ADDR_WIDTH > $clog2(BRAM_DEPTH)) begin
            $warning("Address width exceeds BRAM depth, may cause issues.");
        end
    end

    logic [12:0] addra;
    logic [12:0] addrb;
    
    always_ff @(posedge clk) begin
        if (!rst_n) begin
            addra <= 'd0;
            addrb <= 'd1;
        end 
        else if (in_valid) begin
            if (addra >= LATENCY - 1) begin
                addra <= 'd0;
            end else begin
                addra <= addra + 'd1;
            end

            if (addrb >= LATENCY - 1) begin
                addrb <= 'd0;
            end else begin
                addrb <= addrb + 'd1;
            end
        end
    end
    
    // 行为级双端口 RAM
    logic [DATA_WIDTH-1:0] ram [0:BRAM_DEPTH-1];
    logic [DATA_WIDTH-1:0] data_out_reg;
    
    // 端口 A: 写
    always_ff @(posedge clk) begin
        if (in_valid) begin
            ram[addra] <= data_in;
        end
    end
    
    // 端口 B: 读
    always_ff @(posedge clk) begin
        data_out_reg <= ram[addrb];
    end
    
    assign data_out = data_out_reg;

endmodule